`timescale 1ns / 1ps

module CG(
    );


endmodule
